`ifndef burst_seq_test_sv
`define burst_seq_test_sv
class hbus_burst_seq_test extends hbus_base_test;
    
    hbus_burst_write burst_write;
    hbus_burst_read burst_read;
    
    hbus_extension ext;
    
    hbus_reg_block hbus_rm;
    
    uvm_reg ctrl_p0;
    uvm_reg ctrl_p1;
    uvm_reg ctrl_p2;
    uvm_reg ctrl_p3;
    
    uvm_status_e status;

    uvm_reg_hw_reset_seq reset_seq;
    uvm_reg_bit_bash_seq bit_bash_seq;
    uvm_reg_access_seq access_seq;

    bit [7:0] value;
    
    `uvm_component_utils(hbus_burst_seq_test)
    
    function new (string name, uvm_component parent);
        super.new(name, parent);
    endfunction
    
    function void build_phase (uvm_phase phase);
        super.build_phase(phase);
        burst_write=hbus_burst_write::type_id::create("burst_write", this);
        burst_read=hbus_burst_read::type_id::create("burst_read", this);
        ext=hbus_extension::type_id::create("ext", this);
        reset_seq=uvm_reg_hw_reset_seq::type_id::create("reset_seq");
        bit_bash_seq=uvm_reg_bit_bash_seq::type_id::create("bit_bash_seq");
        access_seq=uvm_reg_access_seq::type_id::create("access_seq");
    endfunction

    function void end_of_elaboration_phase (uvm_phase phase);
        super.end_of_elaboration_phase(phase);
        uvm_resource_db#(bit)::set({"REG::",env.hbus_rm.get_full_name(),".id_register"},"NO_REG_TESTS", 1, this);
        uvm_resource_db#(bit)::set({"REG::",env.hbus_rm.get_full_name(),".bitwise_and"},"NO_REG_TESTS", 1, this);
    endfunction
    
    function void start_of_simulation_phase (uvm_phase phase);
        super.start_of_simulation_phase(phase);
        hbus_rm=env.hbus_rm;
        ctrl_p0=hbus_rm.ctrl_p0;
        ctrl_p1=hbus_rm.ctrl_p1;
        ctrl_p2=hbus_rm.ctrl_p2;
        ctrl_p3=hbus_rm.ctrl_p3;
    endfunction
    
    task run_phase (uvm_phase phase);
        super.run_phase(phase);
        `uvm_info(get_name(), "Start run phase", UVM_MEDIUM)
        phase.phase_done.set_drain_time(this, 5);
        phase.raise_objection(this);
        
        // burst_write.start(env.agnt_main.seqr);
        // burst_read.start(env.agnt_main.seqr);

        // reset_seq.model=env.hbus_rm;
        // reset_seq.start(null);

        // bit_bash_seq.model=env.hbus_rm;
        // bit_bash_seq.start(null);

        // access_seq.model=env.hbus_rm;
        // access_seq.start(null);

        ctrl_p1.set(4);
        ctrl_p2.set(6);
        ctrl_p3.set(8);
        
        ext.burst_size=4;
        ctrl_p0.write
        (
        .status(status),
        .value(8'h02),
        .path(UVM_FRONTDOOR),
        .extension(ext)
        );

        ctrl_p0.read
        (
        .status(status),
        .value(value),
        .path(UVM_FRONTDOOR),
        .extension(ext)
        );
        
        repeat (2) @ (posedge env.agnt_main.drv.m_hbus_if.clk);
        phase.drop_objection(this);
    endtask
endclass
`endif //burst_seq_test_sv