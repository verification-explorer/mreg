`ifndef hbus_pkg_sv
`define hbus_pkg_sv
package hbus_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import hbus_types_pkg::*;

    // Sequence item
    `include "hbus_extension.svh"
    `include "hbus_seq_item.svh"

    // Components
    `include "hbus_cfg.svh"
    `include "hbus_drv.svh"
    `include "hbus_seqr.svh"
    `include "hbus_mntr.svh"
    `include "hbus_agnt.svh"

    // Sequences
    `include "hbus_seq_list.svh"

    // Adepter
    `include "hbus_reg_adapter.svh"
    `include "hbus_reg_adapter_burst.svh"
endpackage
`endif //hbus_pkg_sv